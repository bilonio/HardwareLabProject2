module main (a,b,rnd,z,status);
input logic [31:0] a,b;
input logic [3:0] rnd;
output logic [31:0] z;
output bit [7:0] status; // could use byte?


endmodule
